module history_buffer(
		clock,
		reset
	);

endmodule