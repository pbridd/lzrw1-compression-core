package topPkg;

`include "fileReader.sv"
`include "string_writer.sv"
`include "driver.sv"
`include "env.sv"
`include "testcase.sv"


endpackage	: topPkg
